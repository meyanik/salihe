/home/myanik/work/teknofest24/alaz/playground/gsclib045/gsclib045/lef/gsclib045_tech.lef